`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:10:07 06/07/2017 
// Design Name: 
// Module Name:    RAM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module RAM(
			  input CLK,
			  input CMWr,  
			  input MRd, 
			  input [31:0]AB, 
			  inout [31:0]MD
    );
	 reg [7:0] mem [0:270000];
	 reg [31:0] count;
	 reg [31:0] _MD;
	 
	 initial count = 32'b00000000000000000000000000000000;
	 initial begin
		mem[32'h00000000] = 8'b00000000;
		mem[32'h00000001] = 8'b00000000;
		mem[32'h00000002] = 8'b00000000;
		mem[32'h00000003] = 8'b00000001;
		mem[32'h00000004] = 8'b00000000;
		mem[32'h00000005] = 8'b00000000;
		mem[32'h00000006] = 8'b00000000;
		mem[32'h00000007] = 8'b00000010;
		mem[32'h00000008] = 8'b00000000;
		mem[32'h00000009] = 8'b00000000;
		mem[32'h0000000A] = 8'b00000000;
		mem[32'h0000000B] = 8'b00000011;
		mem[32'h0000000C] = 8'b00000000;
		mem[32'h0000000D] = 8'b00000000;
		mem[32'h0000000E] = 8'b00000000;
		mem[32'h0000000F] = 8'b00000100;
		
		mem[32'h00000010] = 8'b00000000;
		mem[32'h00000011] = 8'b00000000;
		mem[32'h00000012] = 8'b00000000;
		mem[32'h00000013] = 8'b00000101;
		mem[32'h00000014] = 8'b00000000;
		mem[32'h00000015] = 8'b00000000;
		mem[32'h00000016] = 8'b00000000;
		mem[32'h00000017] = 8'b00000110;
		mem[32'h00000018] = 8'b00000000;
		mem[32'h00000019] = 8'b00000000;
		mem[32'h0000001A] = 8'b00000000;
		mem[32'h0000001B] = 8'b00000111;
		mem[32'h0000001C] = 8'b00000000;
		mem[32'h0000001D] = 8'b00000000;
		mem[32'h0000001E] = 8'b00000000;
		mem[32'h0000001F] = 8'b00001000;
		
		mem[32'h00040020] = 8'b00000000;
		mem[32'h00040021] = 8'b00000000;
		mem[32'h00040022] = 8'b00000000;
		mem[32'h00040023] = 8'b00001001;
		mem[32'h00040024] = 8'b00000000;
		mem[32'h00040025] = 8'b00000000;
		mem[32'h00040026] = 8'b00000000;
		mem[32'h00040027] = 8'b00001010;
		mem[32'h00040028] = 8'b00000000;
		mem[32'h00040029] = 8'b00000000;
		mem[32'h0004002A] = 8'b00000000;
		mem[32'h0004002B] = 8'b00001011;
		mem[32'h0004002C] = 8'b00000000;
		mem[32'h0004002D] = 8'b00000000;
		mem[32'h0004002E] = 8'b00000000;
		mem[32'h0004002F] = 8'b00001100;
		
		mem[32'h00000030] = 8'b00000000;
		mem[32'h00000031] = 8'b00000000;
		mem[32'h00000032] = 8'b00000000;
		mem[32'h00000033] = 8'b00000101;
		mem[32'h00000034] = 8'b00000000;
		mem[32'h00000035] = 8'b00000000;
		mem[32'h00000036] = 8'b00000000;
		mem[32'h00000037] = 8'b00000110;
		mem[32'h00000038] = 8'b00000000;
		mem[32'h00000039] = 8'b00000000;
		mem[32'h0000003A] = 8'b00000000;
		mem[32'h0000003B] = 8'b00000111;
		mem[32'h0000003C] = 8'b00000000;
		mem[32'h0000003D] = 8'b00000000;
		mem[32'h0000003E] = 8'b00000000;
		mem[32'h0000003F] = 8'b00001000;
	 end
	 always @(posedge CLK) begin
		if ( MRd == 0 && CMWr != 1) begin
			_MD[31:24] = mem[AB+ (count<<2)];
			_MD[23:16] = mem[AB+(count<<2)+1];
			_MD[15:8] =  mem[AB+(count<<2)+2];
			_MD[7:0] =   mem[AB+(count<<2)+3];
			count = (count+1) & 32'b00000000000000000000000000000011;
      end 

		else if (CMWr == 1) begin
			_MD = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
			if (count != 0) begin
				mem[AB] = MD[31:24];
				mem[AB+1] = MD[23:16];
				mem[AB+2] = MD[15:8];
				mem[AB+3] = MD[7:0];
			end
			count = count +1;
			if (count == 2) 
				count = 4'b0000;
		end
	end
	
	assign  MD = _MD;
	
endmodule
